
`define DATA_W  32
`define ADDR_W  32
`define WDATA_W  32
`define KNN_ENABLE_W 1
`define KNN_VALID_W 1
`define KNN_LOW_W  16
`define KNN_HIGH_W 16
`define K_NEIGHBOUR 6
`define K_NUM_DATA_PTS 127
`define K_DATA_PTS_INDEX_WIDTH 16
  

