
`define TIMER_WIDTH  64
`define DATA_W  32
`define ADDR_W  32
`define WDATA_W  32
`define TIMER_ENABLE_W 1
`define TIMER_SAMPLE_W 1
`define TIMER_LOW_DW 32
`define TIMER_HIGH_DW 32
  

